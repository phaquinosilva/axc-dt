** 4 bit binary reduced logic comparator

* aproximacao: sem logica do bit 0, logica do bit 1 trocado por a1

* result of a <= b in s3
.subckt comp_approx_4b a0 a1 a2 a3 b0 b1 b2 b3 leq vdd
*DUT
* A xnor B
Xeq3 a3 b3 eq3 vdd xnor

Xb2 b2 nb2 vdd Inv
Xb3 b3 nb3 vdd Inv

Xn3 a3 nb3 n3 vdd nand2
Xn2 a2 nb2 eq3 n2 vdd nand3

Xgreater n3 n2 b1 greater vdd nand3
Xinv greater leq vdd inv
.ends