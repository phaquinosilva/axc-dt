* 8 bit dedicated leq comparator

* default settings
.include params.cir

* subcircuit includes
.include gates/rtl_utils.cir

* non-default includes -- simulation source and comparator version
.include simulation_info.txt

* load
.include load_inputs.cir

* DUT
Xcomparator a0 a1 a2 a3 a4 a5 a6 a7 b0 b1 b2 b3 b4 b5 b6 b7 leq vdut comparator

* output load
Cleq leq gnd 1f

* default energy measures
.measure tran q_dut integ i(Vvdut) from=0n to=2.5n
.measure tran q_in integ i(Vvdd1) from=0n to=2.5n

.tran 0.1ns 2.5n

.end
