** 4 bit binary reduced logic comparator

* aproximacao: sem logica do bit 0, logica do bit 1 trocado por a1

* result of a <= b in s3
.subckt comp_approx_4b a0 a1 a2 a3 b0 b1 b2 b3 leq vdd
*DUT
* A xnor B
*Xeq1 a1 b1 eq1 vdd xnor
*Xeq2 a2 b2 eq2 vdd xnor
Xeq3 a3 b3 eq3 vdd xnor

* not B
*Xa0 b0 nb0 vdd Inv
*Xb1 b1 nb1 vdd Inv
Xb2 b2 nb2 vdd Inv
Xb3 b3 nb3 vdd Inv

* greater
Xn3 a3 nb3 n3 vdd nand2
Xn2 a2 nb2 eq3 n2 vdd nand3
*Xn1 a1 nb1 eq3 eq2 n1 vdd nand4
*Xn0 a0 nb0 eq3 eq2 eq1 n0 vdd nand5

* buf
Xia0 a1 na1 vdd Inv
Xia1 na1 n1 vdd Inv

Xgreater n3 n2 n1 greater vdd nand3
Xinv greater leq vdd inv
.ends